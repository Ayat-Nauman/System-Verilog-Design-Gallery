module FF_memory #(parameter WIDTH = 1024, DEPTH = 512 
)(
input logic clk, rst, read_en, write_en,
input logic [$clog2(DEPTH)-1:0]address,
input logic [WIDTH-1:0]write_data,
output logic [WIDTH-1:0]read_data
);

logic [DEPTH-1:0][WIDTH-1:0]memory; //Linear array - width defines word size, depth defines no of rows

generate
	for(genvar i=0; i<DEPTH ; i++) begin
		always_ff @(posedge clk or negedge rst) begin 
			if(!rst)
			memory[i] <= '0;
			else if(address == i && write_en) // write operation
			memory[i] <= write_data;
		end
	end

endgenerate

always_comb begin
	for(int i=0; i<DEPTH; i++) begin
		if(address == i && read_en)
			read_data = memory[i];
	end
end

endmodule

